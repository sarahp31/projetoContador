library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;    -- Biblioteca IEEE para funções aritméticas

entity ULASomaSub is
    generic ( larguraDados : natural := 8 );
    port (
      entradaA, entradaB:  in STD_LOGIC_VECTOR((larguraDados-1) downto 0);
      seletor:  in STD_LOGIC_VECTOR(1 downto 0);
      saida:    out STD_LOGIC_VECTOR((larguraDados-1) downto 0);
		flag: out std_logic
    );
end entity;

architecture comportamento of ULASomaSub is
   signal soma :      STD_LOGIC_VECTOR((larguraDados-1) downto 0);
   signal subtracao : STD_LOGIC_VECTOR((larguraDados-1) downto 0);
	signal passa : STD_LOGIC_VECTOR((larguraDados-1) downto 0);
	signal saida_intermediaria : STD_LOGIC_VECTOR((larguraDados-1) downto 0);
	signal andi :    STD_LOGIC_VECTOR((larguraDados-1) downto 0);
	
    begin
      soma      <= STD_LOGIC_VECTOR(unsigned(entradaA) + unsigned(entradaB));
      subtracao <= STD_LOGIC_VECTOR(unsigned(entradaA) - unsigned(entradaB));
		andi    <= entradaA and entradaB;
		passa <= entradaB;
      saida_intermediaria <= soma when (seletor = "01") else 
									  subtracao when (seletor = "00") else
									  andi when (seletor = "11") else
									  passa;
									  
		flag <= not(saida_intermediaria(7) or saida_intermediaria(6) or saida_intermediaria(5) or saida_intermediaria(4) or saida_intermediaria(3) or saida_intermediaria(2) or saida_intermediaria(1) or saida_intermediaria(0));
		saida <= saida_intermediaria;
end architecture;